Library IEEE;
Use IEEE.STD_LOGIC_1164.ALL;
entity Compuertas is
	port(
		A : in STD_LOGIC;
		B : in STD_LOGIC;
		S1 : out STD_LOGIC;
		S2 : out STD_LOGIC;
		S3 : out STD_LOGIC;
		S4 : out STD_LOGIC;
		S5 : out STD_LOGIC;
		S6 : out STD_LOGIC;
		S7 : out STD_LOGIC

	);
end Compuertas;